// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CE+AbDZ5C8ch8F2vTqxkJM3t+tg54M2OiyYAZT1wOYs+7tPnzlECOlytznomrbXw
SQZ5/9ahfgQKB4Tnv7Amlc3l5GRxwWgCue71JHqhLrTz6uNYNOprFwi1WhhX7PuR
eaqfxo/Hr/Tg0d9P0hF5EHjLIPHgXGwTBLjN0FbPymI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
hPjVowesIjhGGgttxNSDyBPnNO2NP+OgFC6/4QquP8wMAPobf+tyrfhIxPmMkEa3
Q366mjDQt3XwYRQKiiFJ2D77rJT0MnQfe55XhbeXbyriUe8yni5MBFC8OzuYkZls
zTwSwn/0bnBG02sMpXSokhgigjZ/5PK9mj7bP4SNlM8qVZtBymUhFbuTfbAvTvaY
QeRvdvdlx/9mOGOzZLrc6nS8tl/O8suOOsnIqmJPFEYKXjWDe7h60l1pjAwuH+nX
+IzuQ0Q/fVeeHhB6lPHaQrekvbQkd1PjW7+c29mDHb9M5EeK5/06e3fOVaTPGfuQ
x7w2DFi+cspdMDI+KLSY1NIRqC+XeJ74Zo3N9zxv4CYWiQlEijAWGqfSnKjveFRq
tsi3Xb4dwz9r5OgFR0BI9eATCxAtlZ8PpJNFJmEOVWBxA5nkJheNpFudwp6hWwAd
2IlGW2JvgZjI7h79LaEZejdD6QaqC/RN0Ux1RqCMtolirkvnGBN9ieKZ2vVzpk8G
13dLhWeRn1USDdj6ZkEajbiF6f6Bx3eRv/IjB73NFVyB8l8GVl5Tw6tiDmANAr4q
dGrWwwCzi1jYOmPiS2WMPoyH1OFc9qtHwkzO7VyeLF4xsK8kx9Jda5IA5MccLp1M
aqTXCOVYMW1T7yB7BCIuqzFy3hvx2mPAjMRume+2oEbqWTGrYpwMH8TVveOb10Q/
flWG1E2WrsWW/IY26H0j7/5SwfOY2ousPaw+oAHBRKtnFW9bQMcSrG1DWM3MpQUO
12cDwLwz1z9E9bhGlLLQTT4GLIIEY8TYi4um1NnBkYJWUuv80OAG3uSWnrf+rFoJ
SvwKe2oyGQWwFXr8W4NqbduBn7j+2ubHpC6N8TBVo0l0nC8yzvcRlP+6CNlZWvnQ
p0bVIFxpwHsH/7jMEZxUyylemBkWxk0/hntR1CfvH20E40WBx5pCKLyOvqFO8cQw
KQvSg8Z5ZQXRhV8ilF+KWaV0sA67hXO5aN/0rGa5I4eDEl6HJ0U3Q294xKrERB3O
kcpMDIQXKs3Mokt8kVPRqtz1sf7iJZ2zEb9nLoee62gQD1RZbiToadmSsO7pSxuf
rYSrBlWARWdXYzOo6Il+iBRdm26Tkwf4owWD4KJia7zNEocX+zEi25qGPviAhhzK
GqX2k5MMK9GLbnup/f9Bdrr/l5t0aj+Of1EGOMrHtWeWrtuhO9wy3/SwM5W5KVDs
2FD62HxI9xDx/rFoDJLluQ/IITyBbNrZQkFA9bTNBsziPfAswm7WuVxOpSoi6xrl
KnoXmKQtt0C+AeyVCtFYkjPZmxFeBOQF0BEBY3IAcji+pL0DlQOGUVvHkr4FLWpn
9xcYo3yYEKurtlH2Om03h7YMmZ+iQQ0TODtMZ4Iqfjdj43Tut9R/tOJB8xkWKTd7
GIXP9XabXxWhfwgEUDQZJy+c29PkT0hmLMfC8or8a/7C5rtkIM2nrMHvZ/m+RtlR
qjyrC2bKwIl8ldQs5LdyF5QPlB9ZJsfnLlTD/Kwlz2NvIAt3RWa3t/pssfdTt6Na
U0EmJsqLKJfd6wtffbNdGIkqnv9ZVo5j7xuZJaDkY4ngyAmmbC2HmK8o4Wrj3dI1
U0FOmyaIdS3iG6bc1MmjNkK4SJHFF+4GEz0JWjTRykf6rQqjFEq+5Fm4YDuOzFJj
xY8D7s5As3FGv4/xDwvOPtaBy475aldrPnxxPOygmC/ulDHGV4KvXuqW9xccbCQc
0gVrx4kbLIw5mdxnnhuCLQTetSmUXCJ3znFQHH0YCkrF1bDC7Q108zjySN5k686u
1FHTz9gPbxfHYrtrdDUNiHLt0xtPmbgdT1CcNLig0VL7uduD7ga3cwr+612Jpm/A
tnxFTyFS6N89I2YnleXDxaXix3U4jqLmtHWFNfvtLImLL1MgfXXTnXlTkbpmIRpN
XPMJMs5+YYtu6C0miSZW8h+MGXs2gw2SZk5bVde++Ulm07vL1ujN2qL+fdXsUOPk
IdIgdCWtU8+Au86bgjxemtV00DhjpFXD92HRfUPC8P/BS8xsuzbzzBaKTvqnOBm0
sU9iZ94Vn/yCgl42yujs0YxPoT80fnawtErgG8b4CWGgvo/zrXAl0WB5XHBaBw8z
DyxesXp2rSKjsKR+3umo0aipw5GqNliCRgZxLPrK9052DV7j/bICN5P3e50n9oSW
cfRKavCuKeEEm07IHuy/IU4lLcJcRLDAmFVmQTDUu+QXM2J62MH8PWXWdR6weh3p
dU2RMt81h+NgVqAqlA8d247ZqgRfKeXhkkyWY6eaNnaf8FgTy79Knvu6+R3wEEpn
/zaGsIJcPlnksS/Epzmmc28ouv6rRYVVWMp5C0mHHmg/N6KeHqKyM717AnVyQJhi
PuT99NlUy373Eqd5K4hclfsPSXms0AegnkylJjV7BRFsItJQtde+ZGAMIrJd/jeE
6cjtXcw9gGxdZbWQ5zzRY9domZ1Cdua333Q8u5rx86nRtJb+hrLWFbfCrOPE9PeD
LUOTVA9pCwi8DeW9NjgBoi5d7ytxDPovyyPfQXjkiGYqlZrmE9B4V5aGfhdmkLLW
9FwDrh4vE0AZfuFPVMoEMEIk5HPRhvL8WRFgx0XH1oAUFo8+f8B/MoqiBqWgQs9M
d8pzRvj2N3P5Mtti15085qlUcXqxyy4cHpPDjTPwVumWJYOwrBLqXfStin/V+jRs
9G1ydq2NwXNkk5PSeidXFDe2/jYn3LuZYh1wLPfq4D0OmLonADqbtSuUuZPoilCC
ZMOJ7P5jN5UYU99XaMgcwPBwyniroIB8z1QcnV33hoTFoDYDD5pfqYxZXTO+Pofm
8KRKU48jJyEXMNQklKJSW0D7K0fy5O7gNes08ZN3RpGHheNjRzvvQUfXtyk6D5q0
47aOWyE6/64tAHgEYk5IALWt31HNgklalmSCKv1vP83VItKVX8rqp3fo0gM91O2/
zBxgi5rzpXtXXoNWqH3jJexO3n7JoxjRjEjFocBgPtGLsdpYQDg7hernTa5tKGOb
nsqQ/VQWVjnLbvazHR/0N/pCHzvfRZbnRSCi3D0HF8a2DS/Fm8jH+dTHuHc5RwRI
0hcj/7ADQLQgreR2OlXwdx+MJS2VTUkNDHasyKgv5kUh+0MiIlgyT1aKebKy3L8y
VKLXv5LaTcUg9J5Mlwylme4fARsFG59wa61aUVBefUL+ngBCfywShqHoRSSH59eJ
OLR4uv/w2SfrficrofsgGMMpW4bLRdhZLwEMOGqxOc0zqQ8fJgylHHNqUDUSrl7H
KqljjgES7q/vMp2qSR5gxIW45f/YScSqxe0UIoanb7DTsXwimb3z+hnAksh53PKR
qGBXU424tABA/cusZjhgAPyB9pxsIjq9zbM6Bni0Hu92xLNHHY0FvWz7pdUpX6Fo
eItRnTGSwDTV4DTR2NoJMFXQyevNJSRt3NdlW98iAplKQkr190ivctpvcCM61R+o
X4UqV2MyCyiAYfn0wuTdODBEgXdLCpSlqDEI1Iye0R4ogm4aHk16HDWDnmfjTTiw
Zs57q8C1zpsMJyMUL3yVX7l0PTv6tRfV3uiPf7QTpb7cDynPq1BHL6c256/xqYQp
qk9O7SyDoX8rY+1PAHPZOAX36oUakZBIixeeAYG5K8GAvfy9Sjl7SanJLk0g7E6J
g3CUdaGlP9RGnImQDAbq6GVlLKSpSUCILhgqxCdPBSMdZGIXp4/sHvm7zBemk33D
Lu8VQbgM4hDwJDM3cP0KQPwnvyxk6baaqRCIOnGmDi65fMW/PJDRIetnpU0rEXp/
++ZAloCIPpjWD4yiddc9b4EwxQmwGt41YaiV+vSGUDIc3P+8LBP9LHUAQqgwME1O
MnZQhBjqsnHbJi31T2VzVyJ3zLBAGrvgp169qgh1LSVfWK3BLaI18ra94IMPE+ZV
gnmNsVRaMUj3/GlRjPcnNiUs4Fl+gNTgdFHV2vKRfLaSOL0NwbwVSW5p1lahoiwJ
KHXrfqeE133XYjPSb2gBzulBhDdGiYj69M2iWLqv182jiemmvEtnfoFkf7q6hIAw
/vdBftgeBhl8YApT8/YksH+DNEIztdV1+WO2WVLSKmCC4QQXds3oDqo2WXrIlSH6
zNwBXNuqjbC7iiIt1vdpa1ODnNJ29swbFUcgJfe884ebsyHkUg6xQ+z427e0Q7Ye
UM3aQQ0LYMB/vtyVkWSK1v54LY4sTMoGXrni2DolKPGJzCHlUgM6M3qbZf3eoUxo
kS2lLhxLUPuHF3zAZ5F1KtxaKhM/MNi2gY/EOHyKI+mR3aXKUv9FbfforuWLYflV
5+qFXsVAapKrMpCQPdTI1u5R9V/Y3jxJ8h6zRhFuYDywXwb6y9NhO+lRm/Slbrrt
RdLQvG6HnCLU0sXMoLxuIsqp2WAGa31+7vLZbYMVMg/K/elxQ66oRM0jxUNMhkKt
BwlIP5szJEeWpVtz16ar/oWmjQ5mWkdA3LlpL1GPWw7DNHxyPyCTRN0den5nJ9Vt
34Usm9BuoXoEvkiqvKK9Im57SBxYUomArII9ycHXbo4nde31ajs6REcJ09mAM4fg
RUdRmswu8SA95pPx34Mtc0aCVVGMk8Ok2xcryuP6mp0Z5q+C+u00m3o1mjv9KZAs
TnPDz49OMAbzXGKNxlL7Ck7AfZy39AF+nusB840S3HVxTUdi+Krj0/quC+7oZdPm
/Xu2/EKkOdU1Dw0i4akL9BoYIaMzPjmEActoqSpt6Gy+R9yOtO5wD+6jiLNpyDMB
UNEdXCVC2nZlIcuw0yr6Ni5JEPulUhxvfzEXBi+Jci6AtqxkLbUVkfF109UVWJ5K
9oj4CNtQSnttZv+f3DZBhTs8h1aXW08iBPqc5Fv6lkn685bjwtDdgNWp5lzJUMuH
VWs+zBle4AMHeo2pZCUZBkzm3ZyGRuPMDPPrdwmg1gmAm6CmtLFtGvvtQVU0Hsat
d67BZcm6y/tUBPjrmVvcmtoocEgMU/Sj6CwlbOBeAU1xVoOdCWTnhA3WSjKxfjIR
mCNEuaB87xmnnzUdyZzHjwqCkOzpwveUvNSie0sylLeM11m5bjs1+NYi064esbbl
U7fiPqs7xEqPOX1YOyyAueb7gQGsoFE09v6ihN05loSUJSZbZHV0NhYB1ZI6ZkgX
/Zm/BuVMzzLhTSj+VJlgMK9kRSTcn/wDK7PZBxeDF31KgVtmILq3zkD6m/3EcKwj
PIKlF/MY6lekcWfivoQ2lqQzwBP8k9O4jJyMvLOYrWdC6WqFNcYYM/XuZQcytHHg
rg4pmU9PDK/K49zYuLes0sOgLoWtb/6ujmX5Nmd5t+F2//u1JNeKkTV92suKk6PS
UqIxfXmE5Qoe23TcTQDwY9ynJtLtGp84vPskB9hmrysqdwbc4C1R6HtEfap959nS
54wle9kYm+cXTMkaVgt/lgq/UKh/Om55N+3h7QoGP1VaOXxKvoLu3xjxyL0gU8RT
Ht6jW36tCVujU5mp7062TTZ+45l2xLaEd1Qa6RpYDdrJUoup3L2hfr76Z1yKk80f
WPRHEM0z6a0O+FCIxQDANPmzm2FyVhXm7u/U/DdIZMsa16G2xJ5suNmKjCf1pTsd
UneWJxXCb5WEW3viNsiHIoM8828am7rBL/vIYbX0dDt38OPBS1yCC3BfF5nANtmX
iQRpQrF6WACz8DeVgHYEn+nDTQoMKCq6WIiKxZFw+jVXC7nDNdMKw22TdEWa4nCx
n9wzq3D3OLDHtUa9OQYYb6H9k2NSnQk53MJb2L+ZS3fbREfm2o16Xx89YnLstB60
Uyoa5CJcybQ4rUwc65sU8tiRqwMnSF2k0w0S+ojV5wj/xoG2fW8kuZmdLsxQ7QMx
fD/CWgyssyfvSy2NQH9mNqSBTkal379XEaNyQXGPR16WECMhhVjsX71docZMKdqe
YUScbRKAfSWjkrHJoEEqZfivJ0DwUcYUGq1AbRMkBj82TAqx7DlHc+5cP0L5xmFs
+wzxhrWDsZSzuXK9KzhknAfU/fS5oVuBQ/neM89VnvBFpcgoFMZ63sCQw4paLWan
hcq93fPQky+xUsIlwGvwph9SoVTJvLcoV/aDBUVucRlY0eU0Fkkzm3L0S+FclJtl
wmJscamNieqkkEzWv4I8op+Vx+kOu58USZsHJ93OgdGqFdYICKxkMT1TfTXamIY7
+nuLDFb6LlkdmtcLmtqGDeYEw2ufRAMQes+5ZH64w6cIUQFU6LAOa4gNWmsiQNbW
inYANvoOfAAA/vdqhtKnQYwemaCxxLkApVdYNEI7FRI7+gFky4vZRsUDH+BOyBsU
2z8Ka1a10xEp6WPhZENQe/g8fFnRALDXbObFSpfyTDKHAD5kbu6Oe3NoGLnwh5vq
fF7R2tk9XCerultJgZrXf32F/AC2/hd65O8QYapUziqtQz8vVhaODtNN9eGPxY1m
LHJzrs3/Po3Eb7oLYFhMCghxs5Vh6/LWGSsg+Kksqnb71BhQP1hDGQWEX5vQYy6s
1RuU6li5M6RZoYgc5kq5cOSuy1Kj8lPowMKMqqGifR+Vb6S2zH97eevWs1c6eV2j
gVttX1mZizwnZhupspnUnQxiy+sK6k+yzwUASQhpxyNNTFzPtNPRCTXhb/ML6Eok
zJ1eXK1ozbafKsauNzy3oZlfn5Z2S2DNyA+OYsruz03jMxdDOeiG8gYHmIGb6FYo
QkFvQXykaVuwM7PyLyGDqtvJdHNLscBjryAJk4upSD7coLDo1IzxqfXzIIiEJnGa
Qno23p1PL8reY4KmaXqQB6+Y2kUAKYEW4mcjaR0Ud47v5E2QaYm8LpNwixPbQ5KW
r0VZKSHZnIOwGMqbi6VzXPgB0Ied1pDUUMZpAuiKI7UdSGCWMkCQSFvRzxuiYzWK
6Vqyqy6PRmRKu8QpoWTgKiAiNjnpA5oa7RY+U/FE5rHInRpsb3AK5zmiopS2MzhD
n6XBdEo710rlDL+32uHEvBaiKGEUrEnWHMMHKUHtNBK7nfq+tNhCXvR96TdhL+vD
UliCGlCaG6GH2Uatvvn4iprDPUAEaAvkMwzThp/BCS9ricDkEW81ukyUunWHNJ02
R5+rgwJxToOO68z+y+klg/cRDUx0Y5dH4Hnn/Bnpeb+NnZR7u1RzyqdeG2tSbRQS
r9SLE5JOe7gSwRMHD0xc30U9oz+aYJVM0VUUD0wk/LC4Gw/Vz2Qt6emVPj+xafsN
fJ+mwwE5hTxOagMoLQ+nTObfj273yjupJNdTFFfC8llvtOUuoxIq7spnr9Tdzxot
VZQZoS46aau+qTT9BiFf8KPNgnwLKEj0ttFgqgFJIwvebd/pjS3Sfr4Yyu8FdeIi
u+8uU31f4HrxUa91StH159OTvEQPhrIW/avBi3OxiOZeghMTPAPH5EeJ0IyeJBw9
EOXiuXhH3CTD9E45qAaKKp7CYRv3Yua1b4+ZuXDA3SUEFUsXod/6VGMNMruZPxVX
hZtB1up+/ErntYvTGfg39SLGKBGSorS5lFOMrdPsN3Dr4Z/TbSh4Sq67YVnbFFwj
ISbyFwjo53RkDD+/zG1+EPMQFkZCvXYnuFrKQ45TubKpZpXVpBAiLs57doEHVlsO
J9R4NcU67llKu69PhqW7P/H0srxTVhrQBRAfYAXjmNtkFc3cmVmxDRGWyyKERTN6
GGRyd/p6vSBcTJg5kzwa1A==
`pragma protect end_protected
